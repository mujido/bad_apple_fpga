module SD_Card
(
    input chip_select,
    input clk,

    input miso,
    output mosi,

    input RST
);


endmodule
